`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer:       
// Create Date:    12:26:26 04/10/2012 
// Module Name:    control
// Project Name: 	 Lab2
// Description: 	 
//////////////////////////////////////////////////////////////////////////////////
module control(input wire [5:0] opcode,
					output reg [1:0] WB,
					output reg [2:0] M,
					output reg [3:0] EX);


endmodule
